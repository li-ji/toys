
V_1 1 0
R_2 1 2
R_3 2 3
C_4 2 4
C_5 3 0
E_U 4 0 3 0

.end
