
V_1 v_b v_a 32v
V_2 v_c gnd 20v

R_1 v_a ground 2k
R_2 v_c v_b    2k
R_3 v_b ground 4k

.end
