
V_s 1 0 5V
R_1 1 2 1k
C_1 2 0 10p
E_{oa} 4 0 OpAmp 2 3
R_2 4 3 1k
R_3 3 0 1k

.end
