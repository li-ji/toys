
I_{S1} 0 1
I_{S2} 0 3
I_{S3} 1 3

R_1 1 0
R_2 2 0
L_3 3 0
R_4 1 2
C_5 2 3
C_6 1 3

.end
